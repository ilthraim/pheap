module weird_mux #(parameter LEVELS=4) (
    input logic [$clog2(LEVELS):0] sel, [LEVELS:0] a,
    output logic [LEVELS:0] y [$clog2(LEVELS):0]
);

    

endmodule
